CREATE OR ALTER PROCEDURE UI$BLOCK_PARAM_UPD (
    I_BLOCK VARCHAR(30),
    I_PARAM VARCHAR(30),
    I_PARAM_DIRECTION VARCHAR(30),
    I_DATA_TYPE VARCHAR(30),
    I_ORDER_NUM SMALLINT,
    I_CALL_ORDER_NUM SMALLINT,
    I_GROUP_NAME VARCHAR(100),
    I_CAPTION VARCHAR(100),
    I_ENABLER_PARAM VARCHAR(30),
    I_INDEX_IN_KEY SMALLINT,
    I_INDEX_IN_PARENT SMALLINT,
    I_INDEX_IN_NAME SMALLINT,
    I_VISIBLE SMALLINT,
    I_REQUIRED SMALLINT,
    I_READ_ONLY SMALLINT,
    I_DEFAULT_VALUE VARCHAR(1000))
AS
BEGIN
  UPDATE UI$BLOCK_PARAM T
  SET
    T.PARAM_DIRECTION=:I_PARAM_DIRECTION,
    T.DATA_TYPE=:I_DATA_TYPE,
    T.ORDER_NUM=:I_ORDER_NUM,
    T.CALL_ORDER_NUM=:I_CALL_ORDER_NUM,
    T.GROUP_NAME=:I_GROUP_NAME,
    T.CAPTION=:I_CAPTION,
    T.ENABLER_PARAM=:I_ENABLER_PARAM,
    T.INDEX_IN_KEY=:I_INDEX_IN_KEY,
    T.INDEX_IN_PARENT=:I_INDEX_IN_PARENT,
    T.INDEX_IN_NAME=:I_INDEX_IN_NAME,
    T.VISIBLE=:I_VISIBLE,
    T.REQUIRED=:I_REQUIRED,
    T.READ_ONLY=:I_READ_ONLY,
    T.DEFAULT_VALUE = :I_DEFAULT_VALUE
  WHERE T.BLOCK=:I_BLOCK AND T.PARAM=:I_PARAM AND 1=1;
END