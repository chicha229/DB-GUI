CREATE OR ALTER PROCEDURE UI$BLOCK_REF_BIND_CR (
    I_REF INTEGER,
    I_BLOCK VARCHAR(30),
    I_DESTINATION_PARAM VARCHAR(30))
RETURNS (
    REF INTEGER,
    "BLOCK" VARCHAR(30),
    DESTINATION_PARAM VARCHAR(30),
    SOURCE_PARAM VARCHAR(30))
AS
BEGIN
  FOR
    SELECT R.ID, R.BLOCK, RP.PARAM, B.SOURCE_PARAM
    FROM UI$BLOCK_REF R
    JOIN UI$BLOCK_PARAM RP ON RP."BLOCK" = R.REFS_TO AND RP.PARAM_DIRECTION IN ('IN', 'IN_OUT')
    LEFT JOIN UI$BLOCK_REF_BIND B ON B.REF = :I_REF AND B.DESTINATION_PARAM = RP.PARAM
    WHERE
      R.ID = :I_REF AND
      R."BLOCK" = :I_BLOCK AND
      1=1
    INTO :REF,:BLOCK,:DESTINATION_PARAM,:SOURCE_PARAM
  DO SUSPEND;
END