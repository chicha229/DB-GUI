CREATE OR ALTER PROCEDURE UI$FORM_CHILD_PARAM_CR_D (
    I_FORM_CHILD INTEGER,
    I_PARAM VARCHAR(30))
RETURNS (
    FORM_CHILD INTEGER,
    PARAM VARCHAR(30),
    VISIBLE SMALLINT,
    REQUIRED SMALLINT,
    READ_ONLY SMALLINT,
    SOURCE_CHILD INTEGER,
    SOURCE_PARAM VARCHAR(30),
    AUTO_REFRESH SMALLINT)
AS
BEGIN
  FOR
    SELECT :i_form_child,:i_PARAM,T.VISIBLE,T.REQUIRED,T.READ_ONLY,T.SOURCE_CHILD,T.SOURCE_PARAM,T.AUTO_REFRESH
    FROM UI$FORM_CHILD C
    LEFT JOIN UI$FORM_CHILD_PARAM T ON T.FORM_CHILD = :I_FORM_CHILD AND T.PARAM = :I_PARAM
    WHERE
      C.ID = :I_FORM_CHILD AND
      1=1
    INTO :FORM_CHILD,:PARAM,:VISIBLE,:REQUIRED,:READ_ONLY,:SOURCE_CHILD,:SOURCE_PARAM,:AUTO_REFRESH
  DO SUSPEND;
END