CREATE OR ALTER PROCEDURE UI$BLOCK_PARAM_DEL (
    I_BLOCK VARCHAR(30),
    I_PARAM VARCHAR(30),
    I_PARAM_DIRECTION VARCHAR(30),
    I_DATA_TYPE VARCHAR(30),
    I_ORDER_NUM SMALLINT,
    I_GROUP_NAME VARCHAR(100),
    I_CAPTION VARCHAR(100),
    I_ENABLER_PARAM VARCHAR(30),
    I_SOURCE_BLOCK INTEGER,
    I_SOURCE_PARAM VARCHAR(30),
    I_INDEX_IN_KEY SMALLINT,
    I_INDEX_IN_PARENT SMALLINT,
    I_INDEX_IN_NAME SMALLINT,
    I_VISIBLE SMALLINT,
    I_REQUIRED SMALLINT,
    I_READ_ONLY SMALLINT,
    I_DEFAULT_VALUE VARCHAR(1000))
AS
 BEGIN
  DELETE FROM UI$BLOCK_PARAM T
  WHERE T.BLOCK=:I_BLOCK AND T.PARAM=:I_PARAM AND 1=1;
END