CREATE OR ALTER PROCEDURE UI$BLOCK_PARAM_CR_D (
    I_BLOCK VARCHAR(30),
    I_PARAM VARCHAR(30))
RETURNS (
    "BLOCK" VARCHAR(30),
    PARAM VARCHAR(30),
    PARAM_DIRECTION VARCHAR(30),
    DATA_TYPE VARCHAR(30),
    ORDER_NUM SMALLINT,
    CALL_ORDER_NUM SMALLINT,
    GROUP_NAME VARCHAR(100),
    CAPTION VARCHAR(100),
    ENABLER_PARAM VARCHAR(30),
    INDEX_IN_KEY SMALLINT,
    INDEX_IN_PARENT SMALLINT,
    INDEX_IN_NAME SMALLINT,
    VISIBLE SMALLINT,
    REQUIRED SMALLINT,
    READ_ONLY SMALLINT)
AS
BEGIN
  FOR
    SELECT
      T.BLOCK,T.PARAM,T.PARAM_DIRECTION,T.DATA_TYPE,T.ORDER_NUM,CALL_ORDER_NUM,
      T.GROUP_NAME,T.CAPTION,T.ENABLER_PARAM,
      T.INDEX_IN_KEY,T.INDEX_IN_PARENT,T.INDEX_IN_NAME,
      T.VISIBLE,T.REQUIRED,T.READ_ONLY
    FROM UI$BLOCK_PARAM T 
    WHERE
      T.BLOCK = :I_BLOCK AND
      T.PARAM = :I_PARAM AND
      1=1
    INTO
     :BLOCK,:PARAM,:PARAM_DIRECTION,:DATA_TYPE,:ORDER_NUM,:CALL_ORDER_NUM,
     :GROUP_NAME,:CAPTION,:ENABLER_PARAM,
     :INDEX_IN_KEY,:INDEX_IN_PARENT,:INDEX_IN_NAME,
     :VISIBLE,:REQUIRED,:READ_ONLY
  DO SUSPEND;
END