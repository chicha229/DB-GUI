CREATE OR ALTER PROCEDURE UI$BLOCK_PARAM_CR (
    I_BLOCK VARCHAR(30),
    I_PARAM VARCHAR(30))
RETURNS (
    "BLOCK" VARCHAR(30),
    PARAM VARCHAR(30),
    PARAM_DIRECTION VARCHAR(30),
    DATA_TYPE VARCHAR(30),
    ORDER_NUM SMALLINT,
    GROUP_NAME VARCHAR(100),
    CAPTION VARCHAR(100),
    ENABLER_PARAM VARCHAR(30),
    INDEX_IN_KEY SMALLINT,
    INDEX_IN_PARENT SMALLINT,
    INDEX_IN_NAME SMALLINT,
    VISIBLE SMALLINT,
    REQUIRED SMALLINT,
    READ_ONLY SMALLINT,
    L_BLOCK_NAME VARCHAR(100),
    L_PARAM_DIRECTION_NAME VARCHAR(100),
    L_DATA_TYPE_NAME VARCHAR(100))
AS
BEGIN
  FOR
    SELECT
      T.BLOCK,T.PARAM,T.PARAM_DIRECTION,T.DATA_TYPE,T.ORDER_NUM,T.GROUP_NAME,
      T.CAPTION,T.ENABLER_PARAM,T.INDEX_IN_KEY,T.INDEX_IN_PARENT,T.INDEX_IN_NAME,
      T.VISIBLE,T.REQUIRED,T.READ_ONLY,
      L_2.NAME AS L_BLOCK_NAME,L_4.NAME AS L_PARAM_DIRECTION_NAME,L_5.NAME AS L_DATA_TYPE_NAME
    FROM UI$BLOCK_PARAM T
    LEFT JOIN UI$BLOCK L_2 ON L_2.ID = T.BLOCK
    LEFT JOIN UI$PARAM_DIRECTION L_4 ON L_4.ID = T.PARAM_DIRECTION
    LEFT JOIN UI$DATA_TYPE L_5 ON L_5.ID = T.DATA_TYPE
    WHERE
      (T.BLOCK = :I_BLOCK OR :I_BLOCK IS NULL) AND
      (T.PARAM = :I_PARAM OR :I_PARAM IS NULL) AND
      1=1
    ORDER BY T.BLOCK, T.ORDER_NUM
    INTO :BLOCK,:PARAM,:PARAM_DIRECTION,:DATA_TYPE,:ORDER_NUM,:GROUP_NAME,:CAPTION,:ENABLER_PARAM,:INDEX_IN_KEY,:INDEX_IN_PARENT,:INDEX_IN_NAME,:VISIBLE,:REQUIRED,:READ_ONLY,:L_BLOCK_NAME,:L_PARAM_DIRECTION_NAME,:L_DATA_TYPE_NAME
  DO SUSPEND;
END