CREATE OR ALTER PROCEDURE UI$BLOCK_REF_PARAM_DEL (
    I_REF INTEGER,
    I_BLOCK VARCHAR(30),
    I_PARAM VARCHAR(30),
    I_ORDER_NUM SMALLINT,
    I_IS_MAIN_PARAM SMALLINT)
AS
 BEGIN
  DELETE FROM UI$BLOCK_REF_PARAM T
  WHERE T.REF=:I_REF AND T.BLOCK=:I_BLOCK AND T.PARAM=:I_PARAM AND 1=1;
END