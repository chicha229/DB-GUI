CREATE OR ALTER PROCEDURE UI$CR_BLOCK_REF_PARAM
RETURNS (
    REF INTEGER,
    "BLOCK" D_IDENT,
    REFS_TO D_IDENT,
    PARAM D_IDENT,
    ORDER_NUM SMALLINT,
    IS_MAIN_PARAM D_BOOLEAN)
AS
BEGIN
  FOR
    SELECT
      RP.REF, RP."BLOCK", R.REFS_TO, RP.PARAM, RP.ORDER_NUM, RP.IS_MAIN_PARAM
    FROM UI$BLOCK_REF R
    JOIN UI$BLOCK_REF_PARAM RP ON RP.REF = R.ID AND RP."BLOCK" = R."BLOCK"
    ORDER BY R."BLOCK", R.ID, RP.ORDER_NUM
    INTO :REF, :"BLOCK", :REFS_TO, :PARAM, :ORDER_NUM, :IS_MAIN_PARAM
  DO
    SUSPEND;
END