CREATE OR ALTER PROCEDURE UI$FORM_CHILD_REF_BIND_CR (
    I_FORM_CHILD INTEGER)
RETURNS (
    FORM_CHILD INTEGER,
    FORM VARCHAR(30),
    "BLOCK" VARCHAR(30),
    REF INTEGER,
    REF_BLOCK D_IDENT,
    DESTINATION_PARAM VARCHAR(30),
    SOURCE_CHILD INTEGER,
    SOURCE_BLOCK VARCHAR(30),
    SOURCE_PARAM VARCHAR(30))
AS
BEGIN
  FOR
    SELECT C.ID, C.FORM, C."BLOCK", R.ID, R.REFS_TO, DP.PARAM, RB.SOURCE_CHILD, RB.SOURCE_BLOCK, RB.SOURCE_PARAM
    FROM UI$FORM_CHILD C
    JOIN UI$BLOCK_REF R ON R."BLOCK" = C."BLOCK"
    JOIN UI$BLOCK_PARAM DP ON DP."BLOCK" = R.REFS_TO AND DP.PARAM_DIRECTION IN ('in', 'in_out')
    LEFT JOIN UI$FORM_CHILD_REF_BIND RB ON RB.FORM_CHILD = C.ID AND RB.REF = R.ID AND RB.DESTINATION_PARAM = DP.PARAM
    WHERE
      C.ID = :I_FORM_CHILD AND
      1=1
    ORDER BY R.ID, DP.PARAM
    INTO :FORM_CHILD,:FORM,:BLOCK,:REF,:REF_BLOCK,:DESTINATION_PARAM,:SOURCE_CHILD,:SOURCE_BLOCK,:SOURCE_PARAM
  DO SUSPEND;
END