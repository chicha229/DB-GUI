CREATE OR ALTER PROCEDURE UI$BLOCK_REF_PARAM_UPD (
    I_REF INTEGER,
    I_BLOCK VARCHAR(30),
    I_PARAM VARCHAR(30),
    I_ORDER_NUM SMALLINT,
    I_IS_MAIN_PARAM SMALLINT)
AS
BEGIN
  MERGE INTO UI$BLOCK_REF_PARAM T
    USING (SELECT NULL V FROM RDB$DATABASE)
    ON (T.REF = :I_REF AND T."BLOCK" = :I_BLOCK AND T.PARAM = :I_PARAM)
    WHEN MATCHED THEN UPDATE SET
      T.ORDER_NUM = :I_ORDER_NUM,
      T.IS_MAIN_PARAM = :I_IS_MAIN_PARAM
    WHEN NOT MATCHED THEN INSERT (REF,BLOCK,PARAM,ORDER_NUM,IS_MAIN_PARAM)
  VALUES  (:I_REF,:I_BLOCK,:I_PARAM,:I_ORDER_NUM,:I_IS_MAIN_PARAM);
/*
  UPDATE UI$BLOCK_REF_PARAM T
  SET T.ORDER_NUM=:I_ORDER_NUM,T.IS_MAIN_PARAM=:I_IS_MAIN_PARAM
  WHERE T.REF=:I_REF AND T.BLOCK=:I_BLOCK AND T.PARAM=:I_PARAM AND 1=1;
*/
END