CREATE OR ALTER PROCEDURE UI$ACTION_BIND_CR_D (
    I_BLOCK VARCHAR(30),
    I_ACTION VARCHAR(30),
    I_PARAM VARCHAR(30),
    I_DESTINATION_PARAM VARCHAR(30))
RETURNS (
    "BLOCK" VARCHAR(30),
    "ACTION" VARCHAR(30),
    PARAM VARCHAR(30),
    DESTINATION_PARAM VARCHAR(30))
AS
BEGIN
  FOR
    SELECT A.BLOCK,A.ID,T.PARAM,:I_DESTINATION_PARAM
    FROM UI$BLOCK_ACTION A
    LEFT JOIN UI$ACTION_BIND T ON T."BLOCK" = A."BLOCK" AND T.DESTINATION_PARAM = :I_DESTINATION_PARAM AND T.ACTION = :I_ACTION
    WHERE
      A.BLOCK = :I_BLOCK AND
      A.ID = :I_ACTION AND
      1=1
    INTO :BLOCK,:ACTION,:PARAM,:DESTINATION_PARAM
  DO SUSPEND;
END