CREATE OR ALTER PROCEDURE UI$FORM_CHILD_PARAM_UPD (
    I_FORM_CHILD INTEGER,
    I_PARAM VARCHAR(30),
    I_VISIBLE SMALLINT,
    I_REQUIRED SMALLINT,
    I_READ_ONLY SMALLINT,
    I_SOURCE_CHILD INTEGER,
    I_SOURCE_PARAM VARCHAR(30),
    I_AUTO_REFRESH SMALLINT)
AS
  DECLARE VARIABLE L_SOURCE_BLOCK D_IDENT;
  DECLARE VARIABLE L_CHILD_BLOCK D_IDENT;
  DECLARE VARIABLE L_CHILD_FORM D_IDENT;
BEGIN
  SELECT C."BLOCK"
    FROM UI$FORM_CHILD C
    WHERE C.ID = :I_SOURCE_CHILD
    INTO :L_SOURCE_BLOCK;

  SELECT C.FORM, C.BLOCK
    FROM UI$FORM_CHILD C
    WHERE C.ID = :I_FORM_CHILD
    INTO :L_CHILD_FORM, :L_CHILD_BLOCK;

  MERGE INTO UI$FORM_CHILD_PARAM P
    USING (SELECT NULL V FROM RDB$DATABASE)
    ON (P.FORM_CHILD=:I_FORM_CHILD AND P.PARAM=:I_PARAM)
    WHEN MATCHED THEN
      UPDATE SET
        P.VISIBLE=:I_VISIBLE,P.REQUIRED=:I_REQUIRED,P.READ_ONLY=:I_READ_ONLY,
        P.SOURCE_BLOCK = :L_SOURCE_BLOCK,P.SOURCE_CHILD=:I_SOURCE_CHILD,P.SOURCE_PARAM=:I_SOURCE_PARAM,
        P.AUTO_REFRESH=:I_AUTO_REFRESH
    WHEN NOT MATCHED THEN INSERT (
        FORM_CHILD,FORM,BLOCK,PARAM,VISIBLE,
        REQUIRED,READ_ONLY,AUTO_REFRESH,
        SOURCE_BLOCK, SOURCE_CHILD,SOURCE_PARAM)
      VALUES (
        :I_FORM_CHILD,:L_CHILD_FORM, :L_CHILD_BLOCK, :I_PARAM,:I_VISIBLE,
        :I_REQUIRED,:I_READ_ONLY,:I_AUTO_REFRESH,
        :L_SOURCE_BLOCK, :I_SOURCE_CHILD,:I_SOURCE_PARAM
      );
END