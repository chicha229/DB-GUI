CREATE OR ALTER PROCEDURE UI$FORM_CHILD_PARAM_CR (
    I_FORM_CHILD INTEGER,
    I_PARAM VARCHAR(30))
RETURNS (
    FORM_CHILD INTEGER,
    FORM D_IDENT,
    "BLOCK" D_IDENT,
    PARAM VARCHAR(30),
    VISIBLE SMALLINT,
    REQUIRED SMALLINT,
    READ_ONLY SMALLINT,
    SOURCE_CHILD INTEGER,
    SOURCE_PARAM VARCHAR(30),
    AUTO_REFRESH SMALLINT,
    L_FORM_CHILD_ID INTEGER,
    L_SOURCE_BLOCK_ID INTEGER)
AS
BEGIN
  FOR
    SELECT :I_FORM_CHILD,P.PARAM,C.FORM, C."BLOCK", T.VISIBLE,T.REQUIRED,T.READ_ONLY,T.SOURCE_CHILD,T.SOURCE_PARAM,T.AUTO_REFRESH,L1.ID AS L_FORM_CHILD_ID,L2.ID AS L_SOURCE_BLOCK_ID
    FROM UI$FORM_CHILD C
    JOIN UI$BLOCK_PARAM P ON P.BLOCK = C."BLOCK"
    LEFT JOIN UI$FORM_CHILD_PARAM T ON T.FORM_CHILD = :I_FORM_CHILD AND T.param = P.param
    LEFT JOIN UI$FORM_CHILD L1 ON L1.ID=T.FORM_CHILD
    LEFT JOIN UI$FORM_CHILD L2 ON L2.ID=T.SOURCE_CHILD
    WHERE
      C.ID = :I_FORM_CHILD AND
      (T.PARAM = :I_PARAM OR :I_PARAM IS NULL) AND
      1=1
    INTO :FORM_CHILD,:PARAM,:FORM, :BLOCK, :VISIBLE,:REQUIRED,:READ_ONLY,:SOURCE_CHILD,:SOURCE_PARAM,:AUTO_REFRESH,:L_FORM_CHILD_ID,:L_SOURCE_BLOCK_ID
  DO SUSPEND;
END