CREATE OR ALTER PROCEDURE UI$ACTION_BIND_DEL (
    I_BLOCK VARCHAR(30),
    I_ACTION VARCHAR(30),
    I_PARAM VARCHAR(30),
    I_DESTINATION_PARAM VARCHAR(30))
AS
 BEGIN
  DELETE FROM UI$ACTION_BIND T
  WHERE T.BLOCK=:I_BLOCK AND T.ACTION=:I_ACTION AND T.PARAM=:I_PARAM AND 1=1;
END